/******************************************************************
* Description
*	This is a register of 32-bit that corresponds to the PC counter. 
*	This register does not have an enable signal.
* Version:
*	1.0
* Author:
*	Ing: Moreno Kevin and Dong Jorge
* email:
* Date:
*	21/04/2020
******************************************************************/

module Pipe
#(
	parameter N=32
)
(
	input clk,
	input reset,
	input enable,
	input  [N-1:0] DataInput,
	
	
	output reg [N-1:0] DataOutput
);

always@(negedge reset or negedge clk) begin
	if(reset==0)
		DataOutput <= 0;
	else if (enable==1)
		DataOutput<=DataInput;
end

endmodule
//pcreg//